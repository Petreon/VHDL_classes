ENTITY MUX2X1 IS
	PORT(	A,B,C: IN BIT;
		S: OUT BIT);
END MUX2X1;

ARCHITECTURE fluxo OF MUX2X1 IS
BEGIN
    S <= (A AND NOT C) OR (B AND C);
END fluxo;
